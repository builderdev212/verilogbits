`resetall
`timescale 1ns / 1ps
`default_nettype none

module constant_one (
    output wire one
);

    assign one = 1;

endmodule